module Jump_Unit(
    input [31:0] instruction,
    output reg Jump,
    
);